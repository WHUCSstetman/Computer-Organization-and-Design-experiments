
module imme_gen(
    );


endmodule
